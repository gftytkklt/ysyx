`timescale 1ns/1ps

module ysyx_22040750_clint(
    input I_clk,
    input I_rst,
    output [63:0] O_mtime,
    output [63:0] O_mtimecmp
);
endmodule
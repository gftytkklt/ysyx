`timescale 1ns / 1ps

module ysyx_22040750_csr(

);
endmodule
`timescale 1ns / 1ps
module ysyx_22040750_mul_unit(
    input I_sys_clk,
    input I_rst,
    input [64:0] I_mul_op1,
    input [64:0] I_mul_op2,
    input I_mul_valid,
    output [127:0] O_mul_result,
    output O_mul_valid,
    output O_mul_ready
    );
endmodule

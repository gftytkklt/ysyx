`timescale 1ns / 1ps
module ysyx_22040750_foward_unit(
    input [63:0] I_data
);
endmodule
